`timescale 1ns / 1ps

module Zero_1(input wire [7:0] Resultado,
              output wire Zero);

assign Zero = (Resultado == 8'b0);   // Compara si el resultado es cero

endmodule
